CDF       
      x      
   y      @              ;   Bpxy                       
   	P   Btxy                       
   P   Bxy                        
   P   Jpar0                          
   'P   Ni0                        
   1P   Ni_x                    ;P   R0                      ;T   Rpsi                       
   ;X   Rthe                       
   EX   Rxy                        
   OX   Te0                        
   YX   Te_x                    cX   Theta                          
   c\   Ti0                        
   m\   Ti_x                    w\   VE0                        
   w`   Vi0                        
   �`   Vi_x                    �`   Zpsi                       
   �d   Zthe                       
   �d   Zxy                        
   �d   bmag                    �d   bxcvx                          
   �h   bxcvy                          
   �h   bxcvz                          
   �h   dlthe                          
   �h   dpsi                       
   �h   dqdpsi                         
   �h   dx                         
   �h   dy                         
   �h   gjy0                    �h   hthe                       
   �l   hthe0                      l   iNixnorm                   p   ixlb2                      t   ixseps1                    x   ixseps2                    |   jNixnorm                   �   	jyseps1_1                      �   	jyseps1_2                      �   	jyseps2_1                      �   	jyseps2_2                      �   kappaN                         
  �   kappaTe                        
  �   kappaTi                        
  �   kappaV                         
  !�   kappa_g1                       
  +�   kappa_g2                       
  5�   kappa_n                        
  ?�   nx                     I�   ny                     I�   phi0                       
  I�   psixy                          
  S�   q_safe                         
  ]�   qinty                          
  g�   sibdryg                    q�   simagxg                    q�   sinty                          
  q�   x_array                      ( {�=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?��W?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�6(?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�V�?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?�w_?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2?��2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                =ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=ǾT?�bA��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��AĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵAĵA� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� A� AsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAsAE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�AE�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A!�A�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�UA�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?A�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�b?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�1&?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�Q�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?�r�?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��t?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?��9?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7K?�7KA   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A       =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       >"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��<   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  ?���4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g4��g56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez56Ez4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��4��                                                                                                                                                                                                                                                                4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���                                                                                                                                                                                                                                                                56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�56O�4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���                                                                                                                                                                                                                                                                56V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V356V3@�#@�"@�"@� @�@� @�$@�#@�"@�"@�!@� @� @�@�@�@�@�@�@�@�@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@�@�,@�,@�+@�*@�*@�)@�(@�(@�'@�&@�&@�%@�$@�$@�#@�#@�"@�!@�!@� @�@�@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@��@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@��@��@��@��@��@��@�� @�� @���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@�]2@�]1@�]1@�]/@�],@�]/@�]3@�]2@�]1@�]1@�]0@�]/@�]/@�].@�].@�]-@�],@�],@�]+@�]*@�]@�]
@�]	@�]	@�]@�]@�]@�]@�]@�]@�]@�]@�]@�]@�]@�]@�]@�]@�] @�\�@�\�@�]@�]:@�]:@�]9@�]8@�]8@�]7@�]7@�]7@�]6@�]5@�]5@�]4@�]3@�]3@�]2@�]2@�]1@�]0@�]0@�]/@�].@�].@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�&@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�%�@�&@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@�&5@��'@��%@��%@��"@��@��!@��#@��"@��!@��@��@��@��@��@��@��@��@��@��@��@��@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@��@��@��@��@��@��@��	@��@��@��@��@��@��@��@���@���@���@���@���@���@���@���@�Ҝ@�қ@�қ@�ҙ@�Җ@�ҙ@�ҝ@�Ҝ@�қ@�қ@�Қ@�ҙ@�ҙ@�Ҙ@�Ҙ@�җ@�Җ@�Җ@�ҕ@�Ҕ@�҅@��t@��s@��s@��r@��r@��r@��q@��p@��p@��o@��n@��n@��m@��m@��l@��k@��k@��j@��i@��i@�҇@�Ҥ@�Ҥ@�ң@�Ң@�Ң@�ҡ@�ҡ@�ҡ@�Ҡ@�ҟ@�ҟ@�Ҟ@�ҝ@�ҝ@�Ҝ@�Ҝ@�қ@�Қ@�Қ@�ҙ@�Ҙ@�Ҙ@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z@�z
@�z@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�z@�z@�z@�z@�z@�z@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y�@�y��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������դ�գ�գ�ՠ�՝�՟�ա�ՠ�՟�՞�՝�՛�՛�՚�՘�՗�Ֆ�Օ�Ք�Փ�Ն��x��x��w��u��t��s��r��q��p��o��m��m��l��j��i��i��h��g��e��e��|�Փ�Փ�Ց�Ր�Տ�Վ�Ռ�Ռ�Ջ�Չ�Ո�Շ�Ն�Յ�Մ�Ճ�Ձ�Հ�Հ��~��~��|�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������f2�f2�f2�f0�f.�f0�f3�f2�f2�f2�f1�f0�f0�f/�f/�f/�f.�f.�f-�f,�f �f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f
�f
�f"�f9�f9�f8�f7�f7�f6�f6�f6�f6�f5�f5�f4�f3�f3�f2�f2�f2�f1�f1�f0�f/�f/�9�9�9�9�9�9�9"�9"�9"�9"�9"�9"�9"�9"�9"�9"�9"�9"�9"�9"�9�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9	�9"�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�9:�D�C�C�A�>�@�A�A�@�>�>�=�<�;�9�9�7�6�5�4�'���������������
�	������4�3�1�1�/�.�-�,�+�*�)�(�'�&�%�$�"�!�!�������������}����������������������~��}��}��|��{��o��b��a��a��`��`��`��`��_��_��^��]��]��\��\��\��[��[��Z��Y��Y��q����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�ѱ8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�o8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�=,8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8�r�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8Ҩ�8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8��h8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8� 8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8�I�8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8��8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`8ӵ`�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :   :                                                                                                                                                                                                                                                                   :�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��    >"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��       "            ����           ?BB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pBB�pB9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B9Z8B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B0#0B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B'a8B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B�B&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB&pB��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B~�B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��B��A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@A�/@<�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   <   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  ;�  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  7@  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  6�  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   AFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AA~AAT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_AT_A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44A44AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A�}A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��A��   
   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E8Q�E9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9gY9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9�<@9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9��B9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�9�u�:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:�K:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:*�s:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:EXT:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:_��:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;:z8;?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�?˷�    >  >� >� ?  ?H ?p ?� ?� ?� ?� ?� ?� @ @ @ @  @* @4 @> @H @R @\ @f @p @z @� @� @� @�  @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� A A� A A	�A A�A  A�A A�A A�    >  >� >� ?  ?H ?p ?� ?� ?� ?� ?� ?� @ @ @ @  @* @4 @> @H @R @\ @f @p @z @� @� @� @�  @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� A A� A A	�A A�A  A�A A�A A�    >   >�  >�  ?   ?H  ?p  ?�  ?�  ?�  ?�  ?� ?�  @  @  @  @   @*  @4  @>  @H  @R @\ @e��@p  @z  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� @�  @� @�  @���@�  @�  @� @�  @� A  A� A  A	� A  A� A  A� A  A� A  A�     >   >�  >�  ?   ?H  ?p  ?�  ?�  ?�  ?�  ?� ?�  @  @  @  @   @*  @4  @>  @H  @R @\ @e��@p  @z  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� @�  @� @�  @���@�  @�  @� @�  @� A  A� A  A	� A  A� A  A� A  A� A  A�     >   >�  >�  ?   ?H  ?p  ?�  ?�  ?�  ?�  ?� ?�  @  @  @  @   @*  @4  @>  @H  @R @\ @e��@p  @z  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� @�  @� @�  @���@�  @�  @� @�  @� A  A� A  A	� A  A� A  A� A  A� A  A�     >   >�  >�  ?   ?H  ?p  ?�  ?�  ?�  ?�  ?� ?�  @  @  @  @   @*  @4  @>  @H  @R @\ @e��@p  @z  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� @�  @� @�  @���@�  @�  @� @�  @� A  A� A  A	� A  A� A  A� A  A� A  A�     >   >�  >�  ?   ?H  ?p  ?�  ?�  ?�  ?�  ?� ?�  @  @  @  @   @*  @4  @>  @H  @R @\ @e��@p  @z  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� @�  @� @�  @���@�  @�  @� @�  @� A  A� A  A	� A  A� A  A� A  A� A  A�     >  >� >� ?  ?H ?p ?� ?� ?� ?� ?� ?� @ @ @ @  @* @4 @> @H @R @\ @f @p @z @� @� @� @�  @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� A A� A A	�A A�A  A�A A�A A�    >  >� >� ?  ?H ?p ?� ?� ?� ?� ?� ?� @ @ @ @  @* @4 @> @H @R @\ @f @p @z @� @� @� @�  @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� @� A A� A A	�A A�A  A�A A�A A�    >   >�  >�  ?   ?H  ?p  ?�  ?�  ?�  ?�  ?� ?�  @  @  @  @   @*  @4  @>  @H  @R @\ @e��@p  @z  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @�  @� @�  @� @�  @���@�  @�  @� @�  @� A  A� A  A	� A  A� A  A� A  A� A  A� ?�          �I۹�ۺ��Iۺ{SҺ��亯���ۺ�1ֺ�Sһ
:���#\�/��<~ݻIۻU�ٻb1ֻn�Ի{Sһ��h��:绐�e���仝c��\⻩�a���໶6^��~ݻ��\��ۻ�XZ�ՠٻ��X��1ֻ�zU���Ի�S��SҼ �(��h���
:�_&��e�������$�c� 8��#\�&�!�)�a�,ɠ�/��3�66^�9Z��<~ݼ?��B�\�E�                                                                                                                                                                                                                                                                    �I۹�ۺ��Iۺ{SҺ��亯���ۺ�1ֺ�Sһ
:���#\�/��<~ݻIۻU�ٻb1ֻn�Ի{Sһ��h��:绐�e���仝c��\⻩�a���໶6^��~ݻ��\��ۻ�XZ�ՠٻ��X��1ֻ�zU���Ի�S��SҼ �(��h���
:�_&��e�������$�c� 8��#\�&�!�)�a�,ɠ�/��3�66^�9Z��<~ݼ?��B�\�E�    8��9I�9���9��9�S�:��:/��:I�:b1�:{S�:�:�:���:�\�:���:�~�:��:ՠ�:�1�:���:�S�;�h;
:�;�e;��;c;#\�;)�a;/��;66^;<~�;B�\;I�;OXZ;U��;[�X;b1�;hzU;n��;uS;{S�;��(;��h;��;�:�;�_&;��e;���;���;��$;�c;�8�;�\�;��!;��a;�ɠ;���;�;�6^;�Z�;�~�;��;��\;��    ��۹I۹����۹�SҺ��/��Iۺb1ֺ{SҺ�:纖�亣\⺯�ຼ~ݺ�ۺՠٺ�1ֺ��Ժ�Sһ�h�
:��e���c�#\�)�a�/��66^�<~ݻB�\�IۻOXZ�U�ٻ[�X�b1ֻhzU�n�ԻuS�{Sһ��(���h�����:绍_&���e�������仙�$��c��8���\⻦�!���a��ɠ���໳��6^��Z���~ݻ�����\���    8I�8��9��9I�9{S�9���9���9��9�1�9�S�:
:�:��:#\�:/��:<~�:I�:U��:b1�:n��:{S�:��h:�:�:��e:���:�c:�\�:��a:���:�6^:�~�:��\:��:�XZ:ՠ�:��X:�1�:�zU:���:�S:�S�; �(;�h;�;
:�;_&;�e;��;��;�$;c; 8�;#\�;&�!;)�a;,ɠ;/��;3;66^;9Z�;<~�;?�;B�\;E�    8I�8��9��9I�9{S�9���9���9��9�1�9�S�:
:�:��:#\�:/��:<~�:I�:U��:b1�:n��:{S�:��h:�:�:��e:���:�c:�\�:��a:���:�6^:�~�:��\:��:�XZ:ՠ�:��X:�1�:�zU:���:�S:�S�; �(;�h;�;
:�;_&;�e;��;��;�$;c; 8�;#\�;&�!;)�a;,ɠ;/��;3;66^;9Z�;<~�;?�;B�\;E�    8I�8��9��9I�9{S�9���9���9��9�1�9�S�:
:�:��:#\�:/��:<~�:I�:U��:b1�:n��:{S�:��h:�:�:��e:���:�c:�\�:��a:���:�6^:�~�:��\:��:�XZ:ՠ�:��X:�1�:�zU:���:�S:�S�; �(;�h;�;
:�;_&;�e;��;��;�$;c; 8�;#\�;&�!;)�a;,ɠ;/��;3;66^;9Z�;<~�;?�;B�\;E�    8I�8��9��9I�9{S�9���9���9��9�1�9�S�:
:�:��:#\�:/��:<~�:I�:U��:b1�:n��:{S�:��h:�:�:��e:���:�c:�\�:��a:���:�6^:�~�:��\:��:�XZ:ՠ�:��X:�1�:�zU:���:�S:�S�; �(;�h;�;
:�;_&;�e;��;��;�$;c; 8�;#\�;&�!;)�a;,ɠ;/��;3;66^;9Z�;<~�;?�;B�\;E�                                                                                                                                                                                                                                                                :G:ěp;#��;e`;�t�;�9=;���;��{<C�<��