CDF       
      x         y                     :   Bpxy                       �  	$   Btxy                       �  �   Bxy                        �  $   Jpar0                          �  �   Ni0                        �  $   Ni_x                    �   R0                      �   Rpsi                       �  �   Rthe                       �  ,   Rxy                        �  �   Te0                        �  ,   Te_x                    �   Theta                          �  �   Ti0                        �  "0   Ti_x                    $�   VE0                        �  $�   Vi0                        �  '4   Vi_x                    )�   Zpsi                       �  )�   Zthe                       �  ,8   Zxy                        �  .�   bmag                    18   bxcvx                          �  1<   bxcvy                          �  3�   bxcvz                          �  6<   dlthe                          �  8�   dpsi                       �  ;<   dx                         �  =�   dy                         �  @<   gjy0                    B�   hthe                       �  B�   hthe0                       E@   iNixnorm                    ED   ixlb2                       EH   ixseps1                     EL   ixseps2                     EP   jNixnorm                    ET   	jyseps1_1                       EX   	jyseps1_2                       E\   	jyseps2_1                       E`   	jyseps2_2                       Ed   kappaN                         �  Eh   kappaTe                        �  G�   kappaTi                        �  Jh   kappaV                         �  L�   kappa_g1                       �  Oh   kappa_g2                       �  Q�   kappa_n                        �  Th   nx                      V�   ny                      V�   phi0                       �  V�   psixy                          �  Yp   q_safe                         �  [�   qinty                          �  ^p   sibdryg                     `�   simagxg                     `�   sinty                          �  `�   x_array                        cx?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  >�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>��0>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�)�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>�|�>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>��i>�@���>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>�c>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=�,>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�>=(�><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��><��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                @���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@�ff@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@�;d@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���@���BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH  BH      >I�>��?��?I�?{S�?���?���?��?�1�?�S�@
:�@��@#\�@/��@<~�@I�@U��@b1�@n��@{S�@��h@�:�@��e@���@�c@�\�@��a@���@�6^@�~�@��\    >I�>��?��?I�?{S�?���?���?��?�1�?�S�@
:�@��@#\�@/��@<~�@I�@U��@b1�@n��@{S�@��h@�:�@��e@���@�c@�\�@��a@���@�6^@�~�@��\    >I�>��?��?I�?{S�?���?���?��?�1�?�S�@
:�@��@#\�@/��@<~�@I�@U��@b1�@n��@{S�@��h@�:�@��e@���@�c@�\�@��a@���@�6^@�~�@��\    >I�>��?��?I�?{S�?���?���?��?�1�?�S�@
:�@��@#\�@/��@<~�@I�@U��@b1�@n��@{S�@��h@�:�@��e@���@�c@�\�@��a@���@�6^@�~�@��\    >I�>��?��?I�?{S�?���?���?��?�1�?�S�@
:�@��@#\�@/��@<~�@I�@U��@b1�@n��@{S�@��h@�:�@��e@���@�c@�\�@��a@���@�6^@�~�@��\<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       @��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��MB�A�}�A��A��A�W�A���Aѓ�A�1�A�φA�muA�dA��SA�GBA��2A�� A�!A{}�Aj��AY��AI1�A8mtA'�TA�0A!@��@�1�@��T@�!@I1�@!?�!    B�A�}�A��A��A�W�A���Aѓ�A�1�A�φA�muA�dA��SA�GBA��2A�� A�!A{}�Aj��AY��AI1�A8mtA'�TA�0A!@��@�1�@��T@�!@I1�@!?�!    B�A�}�A��A��A�W�A���Aѓ�A�1�A�φA�muA�dA��SA�GBA��2A�� A�!A{}�Aj��AY��AI1�A8mtA'�TA�0A!@��@�1�@��T@�!@I1�@!?�!    B�A�}�A��A��A�W�A���Aѓ�A�1�A�φA�muA�dA��SA�GBA��2A�� A�!A{}�Aj��AY��AI1�A8mtA'�TA�0A!@��@�1�@��T@�!@I1�@!?�!    B�A�}�A��A��A�W�A���Aѓ�A�1�A�φA�muA�dA��SA�GBA��2A�� A�!A{}�Aj��AY��AI1�A8mtA'�TA�0A!@��@�1�@��T@�!@I1�@!?�!    ?�                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �e��e��e��e��e��e��e��e��e��e��e��e��e��e��e��e�    �e��e��e��e��e��e��e��e��e��e��e��e��e�����e�                                                                4�p�                                                    4�p�    �c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C    �c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C�c�C���3�c�C                                                                4�W�                                                    4�W�    �bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз    �bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз�bз����bз?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�! ?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!=� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =� =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�q =�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�ǀ=�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�" =�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�=�x�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <U  <T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�<T�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�>I�    @��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��:@��D@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��N@��M@��:                 ����         <��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��I<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<��x<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�+-<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<�Z\<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<��¸�  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  2�  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         =�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�=�C�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>o�>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>Wj@>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ>�Ȁ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                >�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     @���@�ff@���@�;d@���