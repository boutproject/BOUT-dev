../test-drift-instability/uedge.grd_std.cdl