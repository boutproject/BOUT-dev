CDF       
      x      
   y      @              ;   Bpxy                       
   	P   Btxy                       
   P   Bxy                        
   P   Jpar0                          
   'P   Ni0                        
   1P   Ni_x                    ;P   R0                      ;T   Rpsi                       
   ;X   Rthe                       
   EX   Rxy                        
   OX   Te0                        
   YX   Te_x                    cX   Theta                          
   c\   Ti0                        
   m\   Ti_x                    w\   VE0                        
   w`   Vi0                        
   �`   Vi_x                    �`   Zpsi                       
   �d   Zthe                       
   �d   Zxy                        
   �d   bmag                    �d   bxcvx                          
   �h   bxcvy                          
   �h   bxcvz                          
   �h   dlthe                          
   �h   dpsi                       
   �h   dqdpsi                         
   �h   dx                         
   �h   dy                         
   �h   gjy0                    �h   hthe                       
   �l   hthe0                      l   iNixnorm                   p   ixlb2                      t   ixseps1                    x   ixseps2                    |   jNixnorm                   �   	jyseps1_1                      �   	jyseps1_2                      �   	jyseps2_1                      �   	jyseps2_2                      �   kappaN                         
  �   kappaTe                        
  �   kappaTi                        
  �   kappaV                         
  !�   kappa_g1                       
  +�   kappa_g2                       
  5�   kappa_n                        
  ?�   nx                     I�   ny                     I�   phi0                       
  I�   psixy                          
  S�   q_safe                         
  ]�   qinty                          
  g�   sibdryg                    q�   simagxg                    q�   sinty                          
  q�   x_array                      ( {�=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�1?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?�x?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?�L?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?�!?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?��R?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?��]?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?���?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��%?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h?��h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                =ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=ǾT=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=� }=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��F=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��E=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��z=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=��C=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=��_=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=~�a=ǾTA ?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?�s?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?�l?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A $A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A 
=A VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA VA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA nA �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A �A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A "�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A &�A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A   A       =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��    =��>I�>���>��>�S�?��?/��?I�?b1�?{S�?�:�?���?�\�?���?�~�?��?ՠ�?�1�?���?�S�@�h@
:�@�e@��@c@#\�@)�a@/��@66^@<~�@B�\@I�@OXZ@U��@[�X@b1�@hzU@n��@uS@{S�@��(@��h@��@�:�@�_&@��e@���@���@��$@�c@�8�@�\�@��!@��a@�ɠ@���@�@�6^@�Z�@�~�@��@��\@��<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
<#�
�   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       >"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��<   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  <   <�  =   =`  =�  =�  =�  =�  >  >  >(  >8  >H  >X  >h  >x  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  >�  ?  ?  ?
  ?  ?  ?  ?  ?  ?"  ?&  ?*  ?.  ?2  ?6  ?:  ?>  ?B  ?F  ?J  ?N  ?R  ?V  ?Z  ?^  ?b  ?f  ?j  ?n  ?r  ?v  ?z  ?~  ?��6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6SSp6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6��$6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6SS�6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6S �6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6ST�6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6S!(6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6��6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6SUL6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6��l6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�6SU�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?F�?+m?+k?+l?+j?+g?+j?+m?+l?+k?+j?+j?+i?+h?+g?+g?+g?+f?+e?+d?+c?+V?+J?+I?+H?+H?+G?+F?+E?+E?+E?+D?+C?+B?+A?+A?+@?+@?+??+>?+>?+=?+U?+m?+l?+l?+k?+j?+j?+i?+h?+g?+g?+g?+f?+e?+d?+c?+c?+b?+b?+a?+`?+`?+_?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?V�?g�?g�?g�?g�?g?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g?g~?g~?gq?gd?gd?gc?gb?gb?gb?ga?ga?g`?g_?g_?g^?g^?g^?g]?g]?g\?g[?g[?g[?gs?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?g�?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?N�?O?O ?O ?O ?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?O?`?`?`?`?`?`?`?`?`?`?`?`?`?`?`?`?`?`?` ?` ?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?_�?`?`?`?`?`?`
?`
?`	?`	?`	?`?`?`?`?`?`?`?`?`?`?`?`?�B?�@?�A?�??�=?�??�B?�A?�@?�@?�??�>?�=?�=?�=?�<?�;?�:?�9?�9?�,?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�*?�B?�A?�A?�@?�@?�??�>?�=?�=?�=?�<?�;?�:?�9?�9?�8?�7?�7?�6?�6?�5?�4?D?D?D?D?D?D?D?D?D?D?D?D?D?D?D?D?D?D?D?D ?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?C�?D?D?D?D?D?D?D
?D
?D	?D?D?D?D?D?D?D?D?D?D?D?D?D?)?)?)?)?)	?)?)?)?)?)?)?)?)
?)	?)	?)?)?)?)?)?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?(�?)?)?)?)?)?)?)?)
?)	?)	?)?)?)?)?)?)?)?)?)?)?)?) ?<??<>?<>?<=?<:?<=?<@?<??<>?<>?<>?<=?<=?<<?<<?<;?<:?<:?<:?<9?<-?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<?<.?<F?<F?<E?<D?<D?<D?<C?<C?<B?<A?<A?<A?<@?<@?<??<??<>?<>?<>?<=?<<?<<�Ǯ.�Ǯ.�Ǯ.�Ǯ,�Ǯ)�Ǯ,�Ǯ0�Ǯ.�Ǯ.�Ǯ.�Ǯ-�Ǯ,�Ǯ,�Ǯ*�Ǯ*�Ǯ*�Ǯ)�Ǯ)�Ǯ(�Ǯ'�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ�Ǯ �ǭ��ǭ��ǭ��ǭ��ǭ��ǭ��ǭ��ǭ��ǭ��ǭ��Ǯ�Ǯ7�Ǯ7�Ǯ7�Ǯ6�Ǯ6�Ǯ5�Ǯ3�Ǯ3�Ǯ3�Ǯ2�Ǯ2�Ǯ1�Ǯ0�Ǯ0�Ǯ.�Ǯ.�Ǯ.�Ǯ-�Ǯ-�Ǯ,�Ǯ*�Ǯ*�ǋ�ǋ�ǋ�ǋ�ǋ	�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ
�ǋ	�ǋ	�ǋ	�ǋ�ǋ�ǋ�ǋ�Ǌ�Ǌ�Ǌ�Ǌ�Ǌ�Ǌ�Ǌ߽Ǌ޽Ǌ޽Ǌ޽ǊܽǊ۽ǊڽǊٽǊٽǊ׽Ǌ׽ǊֽǊսǊսǊԽǊ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ
�ǋ	�ǋ	�ǋ	�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ�ǋ �ǋ �Ǌ����ܽ��۽��۽��ڽ��ֽ��ڽ��ݽ��ܽ��۽��۽��ڽ��ڽ��ڽ��ؽ��ؽ��׽��ֽ��ֽ��ֽ��Խ��Ľ�³��³��³��²��±��±��¯��®��®��®��­��­��¬��¬��ª��ª��ª��©��¨��¨���ƽ�����������������������������߽��߽��߽��ݽ��ݽ��ܽ��ܽ��۽��ڽ��ڽ��ڽ��ؽ��ؽ��"��� ���"������������"���"���"��� ��� ������������������������������
���������������������������������������������������������������������������+���)���)���)���(���'���'���&���&���&���$���$���#���"���"���"��� ��� �������������Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹy�Ǹx�Ǹx�Ǹv�Ǹu�Ǹu�Ǹu�Ǹt�Ǹt�Ǹs�Ǹq�Ǹq�Ǹp�Ǹp�Ǹp�Ǹo�Ǹo�Ǹn�Ǹl�Ǹl�Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ��Ǹ����J���I���J���G���D���H���J���J���J���I���I���H���G���G���E���E���E���D���C���C���2���"���"��� ������������������������������������������������������5���S���S���R���R���Q���O���O���N���N���N���M���M���L���J���J���J���I���I���H���G���G���E��4/��4-��4.��4+��4)��4+��4/��4.��4-��4-��4+��4*��4)��4)��4)��4(��4&��4%��4$��4$��4��4��4��4��4 ��3���3���3���3���3���3���3���3���3���3���3���3���3���3���3��3��4��4/��4.��4.��4-��4-��4+��4*��4)��4)��4)��4(��4&��4%��4$��4$��4#��4!��4!��4 ��4 ��4��4�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�ǩ��ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ�ǩ��Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�Ǫ�ǇO�ǇM�ǇO�ǇK�ǇH�ǇK�ǇO�ǇO�ǇM�ǇL�ǇK�ǇK�ǇI�ǇH�ǇH�ǇG�ǇF�ǇF�ǇD�ǇC�Ǉ3�Ǉ#�Ǉ"�Ǉ!�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ�Ǉ0�ǇO�ǇO�ǇO�ǇM�ǇL�ǇK�ǇK�ǇI�ǇH�ǇH�ǇG�ǇF�ǇF�ǇD�ǇC�ǇB�ǇB�ǇB�ǇA�Ǉ?�Ǉ>�Ǉ=�ǟ�ǟ�ǟ�ǟ߽ǟܽǟ߽ǟ�ǟ�ǟ�ǟ�ǟ�ǟ߽ǟ߽ǟ޽ǟ޽ǟݽǟܽǟܽǟܽǟڽǟ˽ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ��ǟ̽ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ�ǟ߽ǟ޽ǟ�<�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  <�  :��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:�Y:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�!�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�$�:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�(L:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�+�:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�/:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p:�2p8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  8@  7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7�  7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   7   �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  :�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�H:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Q:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�Z:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�b:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�j:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�s:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:�|:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��:��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��    >"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��       "            ����           ?@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�z�@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�90@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@�R�@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@��@s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @s @g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@g'�@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@[�@@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@Q�@F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� @F� �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  :�  �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  �@  5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   5   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  =��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=��O=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=�yJ=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=��=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=���=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=˘,=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=ˬ�=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=��|=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=˗�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�=�n�   
   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                :::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6:ğ6;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;#� ;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;ejW;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�} ;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;�E�;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��;��<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<R�<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��>"��    <�  =   =@  =�  =�  =�  =�  >   >  >   >0  >@  >P  >`  >o��>�  >�  >�  >�  >�  >�  >�  >���>�  >�  >�  >�  >�  >���>���>�  ?   ?  ?  ?  ?  ?  ?  ?  ?   ?#��?(  ?,  ?0  ?4  ?7��?<  ?@  ?D  ?H  ?L  ?P  ?S��?X  ?\  ?`  ?d  ?g��?l  ?o��?t  ?x  ?|      <� =  =@ =� =� =� =� >  > >  >0 >@ >P >` >p >� >� >� >� >� >� >� >� >� >� >� >� >� >� >� >� ?  ? ? ? ? ? ? ? ?  ?$ ?( ?, ?0 ?4 ?8 ?< ?@ ?D ?H ?L ?P ?T ?X ?\ ?` ?d ?h ?l ?p ?t ?x ?|     <� =  =@ =� =� =� =� >  > >  >0 >@ >P >` >p >� >� >� >� >� >� >� >�  >� >� >� >� >� >� >� >� ?  ? ? ? ? ? ? ? ?  ?$  ?( ?, ?0 ?4 ?8  ?< ?@ ?D ?H ?L ?P ?T ?X ?\ ?` ?d ?h ?l ?p ?t ?x ?|     <� =  =@ =� =� =� =� >  > >  >0 >@ >P >` >p >� >� >� >� >� >� >� >�  >� >� >� >� >� >� >� >� ?  ? ? ? ? ? ? ? ?  ?$  ?( ?, ?0 ?4 ?8  ?< ?@ ?D ?H ?L ?P ?T ?X ?\ ?` ?d ?h ?l ?p ?t ?x ?|     <�  =   =@  =�  =�  =�  =�  >   >  >   >0  >@  >P  >`  >o��>�  >�  >�  >�  >�  >�  >�  >���>�  >�  >�  >�  >�  >���>���>�  ?   ?  ?  ?  ?  ?  ?  ?  ?   ?#��?(  ?,  ?0  ?4  ?7��?<  ?@  ?D  ?H  ?L  ?P  ?S��?X  ?\  ?`  ?d  ?g��?l  ?o��?t  ?x  ?|      <�  =   =@  =�  =�  =�  =�  >   >  >   >0  >@  >P  >`  >o��>�  >�  >�  >�  >�  >�  >�  >���>�  >�  >�  >�  >�  >���>���>�  ?   ?  ?  ?  ?  ?  ?  ?  ?   ?#��?(  ?,  ?0  ?4  ?7��?<  ?@  ?D  ?H  ?L  ?P  ?S��?X  ?\  ?`  ?d  ?g��?l  ?o��?t  ?x  ?|      <� =  =@ =� =� =� =� >  > >  >0 >@ >P >` >p >� >� >� >� >� >� >� >� >� >� >� >� >� >� >� >� ?  ? ? ? ? ? ? ? ?  ?$ ?( ?, ?0 ?4 ?8 ?< ?@ ?D ?H ?L ?P ?T ?X ?\ ?` ?d ?h ?l ?p ?t ?x ?|     <�  =   =@  =�  =�  =�  =�  >   >  >   >0  >@  >P  >`  >o��>�  >�  >�  >�  >�  >�  >�  >���>�  >�  >�  >�  >�  >���>���>�  ?   ?  ?  ?  ?  ?  ?  ?  ?   ?#��?(  ?,  ?0  ?4  ?7��?<  ?@  ?D  ?H  ?L  ?P  ?S��?X  ?\  ?`  ?d  ?g��?l  ?o��?t  ?x  ?|      <� =  =@ =� =� =� =� >  > >  >0 >@ >P >` >p >� >� >� >� >� >� >� >�  >� >� >� >� >� >� >� >� ?  ? ? ? ? ? ? ? ?  ?$  ?( ?, ?0 ?4 ?8  ?< ?@ ?D ?H ?L ?P ?T ?X ?\ ?` ?d ?h ?l ?p ?t ?x ?|     <� =  =@ =� =� =� =� >  > >  >0 >@ >P >` >p >� >� >� >� >� >� >� >�  >� >� >� >� >� >� >� >� ?  ? ? ? ? ? ? ? ?  ?$  ?( ?, ?0 ?4 ?8  ?< ?@ ?D ?H ?L ?P ?T ?X ?\ ?` ?d ?h ?l ?p ?t ?x ?| ?�          6���7��7b1�7���7�~�7�1�8�h8��8)�`8<~�8OXZ8b1�8uS8��h8�_&8���8�8�8��`8�8�~�8��8�XZ8��8�1�8랔8�S8�x9�h9��9_&9�9��9�D9 8�9$�9)�`9.[�9397�~9<~�9A5<9E�9J��9OXZ9T�9X�9]{x9b1�9f�69k��9pT�9uS9y��9~x9��89��h9�M�9���9��9�_&9��V9��9�p�    5I�5��6��6I�6{S�6���6���6��6�1�6�S�7
:�7��7#\�7/��7<~�7I�7U��7b1�7n��7{S�7��h7�:�7��e7���7�c7�\�7��a7���7�6^7�~�7��\7��7�XZ7ՠ�7��X7�1�7�zU7���7�S7�S�8 �(8�h8�8
:�8_&8�e8��8��8�$8c8 8�8#\�8&�!8)�a8,ɠ8/��83866^89Z�8<~�8?�8B�\8E�    �I۵�۶��I۶{SҶ��䶯���۶�1ֶ�Sҷ
:���#\�/��<~ݷI۷U�ٷb1ַn�Է{Sҷ��h��:緐�e���䷝c��\ⷩ�a���෶6^��~ݷ��\��۷�XZ�ՠٷ��X��1ַ�zU���Է�S��SҸ �(��h���
:�_&��e�������$�c� 8��#\�&�!�)�a�,ɠ�/��3�66^�9Z��<~ݸ?��B�\�E�    �I۵�۶��I۶{SҶ��䶯���۶�1ֶ�Sҷ
:���#\�/��<~ݷI۷U�ٷb1ַn�Է{Sҷ��h��:緐�e���䷝c��\ⷩ�a���෶6^��~ݷ��\��۷�XZ�ՠٷ��X��1ַ�zU���Է�S��SҸ �(��h���
:�_&��e�������$�c� 8��#\�&�!�)�a�,ɠ�/��3�66^�9Z��<~ݸ?��B�\�E�    ��۶I۶����۶�Sҷ��/��I۷b1ַ{Sҷ�:緖�䷣\ⷯ�෼~ݷ�۷ՠٷ�1ַ��Է�SҸ�h�
:��e���c�#\�)�a�/��66^�<~ݸB�\�I۸OXZ�U�ٸ[�X�b1ָhzU�n�ԸuS�{SҸ��(���h�����:縍_&���e�������丙�$��c��8���\⸦�!���a��ɠ���ำ��6^��Z���~ݸ�����\���    5��6I�6���6��6�S�7��7/��7I�7b1�7{S�7�:�7���7�\�7���7�~�7��7ՠ�7�1�7���7�S�8�h8
:�8�e8��8c8#\�8)�a8/��866^8<~�8B�\8I�8OXZ8U��8[�X8b1�8hzU8n��8uS8{S�8��(8��h8��8�:�8�_&8��e8���8���8��$8�c8�8�8�\�8��!8��a8�ɠ8���8�8�6^8�Z�8�~�8��8��\8��    5I�5��6��6I�6{S�6���6���6��6�1�6�S�7
:�7��7#\�7/��7<~�7I�7U��7b1�7n��7{S�7��h7�:�7��e7���7�c7�\�7��a7���7�6^7�~�7��\7��7�XZ7ՠ�7��X7�1�7�zU7���7�S7�S�8 �(8�h8�8
:�8_&8�e8��8��8�$8c8 8�8#\�8&�!8)�a8,ɠ8/��83866^89Z�8<~�8?�8B�\8E�    �I۵�۶��I۶{SҶ��䶯���۶�1ֶ�Sҷ
:���#\�/��<~ݷI۷U�ٷb1ַn�Է{Sҷ��h��:緐�e���䷝c��\ⷩ�a���෶6^��~ݷ��\��۷�XZ�ՠٷ��X��1ַ�zU���Է�S��SҸ �(��h���
:�_&��e�������$�c� 8��#\�&�!�)�a�,ɠ�/��3�66^�9Z��<~ݸ?��B�\�E�    5I�5��6��6I�6{S�6���6���6��6�1�6�S�7
:�7��7#\�7/��7<~�7I�7U��7b1�7n��7{S�7��h7�:�7��e7���7�c7�\�7��a7���7�6^7�~�7��\7��7�XZ7ՠ�7��X7�1�7�zU7���7�S7�S�8 �(8�h8�8
:�8_&8�e8��8��8�$8c8 8�8#\�8&�!8)�a8,ɠ8/��83866^89Z�8<~�8?�8B�\8E�    ������b1ַ��䷼~޷�1ָ�h���)�`�<~޸OXZ�b1ָuS���h��_&���丠8����`����~޸�뜸�XZ�����1ָ랔��S��x��h��ƹ_&������D� 8��$��)�`�.[��3�7�~�<~޹A5<�E뜹J���OXZ�T��X��]{x�b1ֹf�6�k���pT��uS�y���~x���8���h��M����ƹ����_&���V�����p�:G:ěp;#��;e`;�t�;�9=;���;��{<C�<��